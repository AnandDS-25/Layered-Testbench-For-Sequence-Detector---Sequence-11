interface intf();
  
  bit clk;
 
  bit [1:0]in;
  bit out;
  int count;
  
endinterface